module simple_clock_vcd(input wire clk);

endmodule
module test();
    initial begin
        $display("hello world");
    end
endmodule
